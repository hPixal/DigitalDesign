library ieee;
use ieee.std_logic_1164.all;

entity Motor is
port(
    med : in std_logic;
    alt : in std_logic
);
end entity;
