library ieee;
use ieee.std_logic_1164.all;

entity Sensor is
port(
    sal_sensor : out std_logic
);
end entity;
