-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Aug 4 2020 16:48:09

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "divider" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

--library ice;
library work;
--use ice.vcomponent_vital.all;
use work.vcomponent_vital.all;

-- Entity of divider
entity divider is
port (
    res_out : out std_logic_vector(7 downto 0);
    rmn_out : out std_logic_vector(7 downto 0);
    den_in : in std_logic_vector(7 downto 0);
    num_in : in std_logic_vector(7 downto 0);
    start_in : in std_logic;
    running_out : out std_logic;
    rst_in_n : in std_logic;
    resultOk_out : out std_logic;
    divZero_out : out std_logic;
    clk_in : in std_logic);
end divider;

-- Architecture of divider
-- View name is \INTERFACE\
architecture \INTERFACE\ of divider is

signal \N__3514\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2527\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2478\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2380\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2328\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2277\ : std_logic;
signal \N__2274\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2259\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2247\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2239\ : std_logic;
signal \N__2236\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2224\ : std_logic;
signal \N__2221\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2214\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2196\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2176\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2170\ : std_logic;
signal \N__2167\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2146\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2139\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2132\ : std_logic;
signal \N__2129\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2107\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2095\ : std_logic;
signal \N__2092\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2080\ : std_logic;
signal \N__2077\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2071\ : std_logic;
signal \N__2068\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2062\ : std_logic;
signal \N__2059\ : std_logic;
signal \N__2056\ : std_logic;
signal \N__2053\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2047\ : std_logic;
signal \N__2044\ : std_logic;
signal \N__2041\ : std_logic;
signal \N__2038\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2032\ : std_logic;
signal \N__2029\ : std_logic;
signal \N__2026\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2017\ : std_logic;
signal \N__2014\ : std_logic;
signal \N__2013\ : std_logic;
signal \N__2012\ : std_logic;
signal \N__2011\ : std_logic;
signal \N__2008\ : std_logic;
signal \N__2005\ : std_logic;
signal \N__2002\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1990\ : std_logic;
signal \N__1987\ : std_logic;
signal \N__1984\ : std_logic;
signal \N__1981\ : std_logic;
signal \N__1980\ : std_logic;
signal \N__1979\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1973\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1960\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1953\ : std_logic;
signal \N__1952\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1946\ : std_logic;
signal \N__1943\ : std_logic;
signal \N__1936\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1930\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1926\ : std_logic;
signal \N__1925\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1916\ : std_logic;
signal \N__1909\ : std_logic;
signal \N__1906\ : std_logic;
signal \N__1903\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1897\ : std_logic;
signal \N__1894\ : std_logic;
signal \N__1891\ : std_logic;
signal \N__1888\ : std_logic;
signal \N__1885\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1870\ : std_logic;
signal \N__1867\ : std_logic;
signal \N__1864\ : std_logic;
signal \N__1861\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1843\ : std_logic;
signal \N__1840\ : std_logic;
signal \N__1837\ : std_logic;
signal \N__1834\ : std_logic;
signal \N__1831\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1825\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1819\ : std_logic;
signal \N__1816\ : std_logic;
signal \N__1813\ : std_logic;
signal \N__1810\ : std_logic;
signal \N__1807\ : std_logic;
signal \N__1804\ : std_logic;
signal \N__1801\ : std_logic;
signal \N__1798\ : std_logic;
signal \N__1795\ : std_logic;
signal \N__1792\ : std_logic;
signal \N__1789\ : std_logic;
signal \N__1786\ : std_logic;
signal \N__1783\ : std_logic;
signal \N__1780\ : std_logic;
signal \N__1777\ : std_logic;
signal \N__1774\ : std_logic;
signal \N__1771\ : std_logic;
signal \N__1768\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1753\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1747\ : std_logic;
signal \N__1744\ : std_logic;
signal \N__1741\ : std_logic;
signal \N__1738\ : std_logic;
signal \N__1735\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1729\ : std_logic;
signal \N__1726\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1720\ : std_logic;
signal \N__1717\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1711\ : std_logic;
signal \N__1708\ : std_logic;
signal \N__1705\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1693\ : std_logic;
signal \N__1690\ : std_logic;
signal \N__1687\ : std_logic;
signal \N__1684\ : std_logic;
signal \N__1681\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1675\ : std_logic;
signal \N__1672\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1666\ : std_logic;
signal \N__1663\ : std_logic;
signal \N__1660\ : std_logic;
signal \N__1657\ : std_logic;
signal \N__1654\ : std_logic;
signal \N__1651\ : std_logic;
signal \N__1648\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1642\ : std_logic;
signal \N__1639\ : std_logic;
signal \N__1636\ : std_logic;
signal \N__1633\ : std_logic;
signal \N__1630\ : std_logic;
signal \N__1627\ : std_logic;
signal \N__1624\ : std_logic;
signal \N__1621\ : std_logic;
signal \N__1618\ : std_logic;
signal \N__1615\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1603\ : std_logic;
signal \N__1600\ : std_logic;
signal \N__1597\ : std_logic;
signal \N__1594\ : std_logic;
signal \N__1591\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1582\ : std_logic;
signal \N__1579\ : std_logic;
signal \N__1576\ : std_logic;
signal \N__1573\ : std_logic;
signal \N__1570\ : std_logic;
signal \N__1567\ : std_logic;
signal \N__1564\ : std_logic;
signal \N__1561\ : std_logic;
signal \N__1558\ : std_logic;
signal \N__1555\ : std_logic;
signal \N__1552\ : std_logic;
signal \N__1549\ : std_logic;
signal \N__1546\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1537\ : std_logic;
signal \N__1534\ : std_logic;
signal \N__1531\ : std_logic;
signal \N__1528\ : std_logic;
signal \N__1525\ : std_logic;
signal \N__1522\ : std_logic;
signal \N__1519\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1504\ : std_logic;
signal \N__1501\ : std_logic;
signal \N__1498\ : std_logic;
signal \N__1495\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1486\ : std_logic;
signal \N__1483\ : std_logic;
signal \N__1480\ : std_logic;
signal \N__1477\ : std_logic;
signal \N__1474\ : std_logic;
signal \N__1471\ : std_logic;
signal \N__1468\ : std_logic;
signal \N__1465\ : std_logic;
signal \N__1462\ : std_logic;
signal \N__1459\ : std_logic;
signal \N__1456\ : std_logic;
signal \N__1453\ : std_logic;
signal \N__1450\ : std_logic;
signal \N__1447\ : std_logic;
signal \N__1444\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal rst_in_n_c : std_logic;
signal rst_in_n_c_i : std_logic;
signal den_in_c_0 : std_logic;
signal den_in_c_5 : std_logic;
signal den_in_c_6 : std_logic;
signal num_in_c_0 : std_logic;
signal num_in_c_1 : std_logic;
signal num_in_c_2 : std_logic;
signal num_in_c_3 : std_logic;
signal num_in_c_4 : std_logic;
signal num_in_c_5 : std_logic;
signal num_in_c_6 : std_logic;
signal rmn_out_c_7 : std_logic;
signal rmn_out_c_3 : std_logic;
signal rmn_out_c_4 : std_logic;
signal rmn_out_c_5 : std_logic;
signal rmn_out_c_6 : std_logic;
signal rmn_out_c_0 : std_logic;
signal rmn_out_c_2 : std_logic;
signal rmn_out_c_1 : std_logic;
signal res_out_c_0 : std_logic;
signal res_out_c_3 : std_logic;
signal res_out_c_7 : std_logic;
signal res_out_c_6 : std_logic;
signal res_out_c_4 : std_logic;
signal res_out_c_2 : std_logic;
signal res_out_c_5 : std_logic;
signal res_out_c_1 : std_logic;
signal den_reg_i_0 : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal load_and_iterate_iterate_reg_1_1 : std_logic;
signal load_and_iterate_iterate_reg_1_cry_0 : std_logic;
signal load_and_iterate_iterate_reg_1_2 : std_logic;
signal load_and_iterate_iterate_reg_1_cry_1 : std_logic;
signal load_and_iterate_iterate_reg_1_3 : std_logic;
signal load_and_iterate_iterate_reg_1_cry_2 : std_logic;
signal load_and_iterate_iterate_reg_1_4 : std_logic;
signal load_and_iterate_iterate_reg_1_cry_3 : std_logic;
signal den_reg_i_5 : std_logic;
signal load_and_iterate_iterate_reg_1_5 : std_logic;
signal load_and_iterate_iterate_reg_1_cry_4 : std_logic;
signal den_reg_i_6 : std_logic;
signal load_and_iterate_iterate_reg_1_6 : std_logic;
signal load_and_iterate_iterate_reg_1_cry_5 : std_logic;
signal num_in_c_7 : std_logic;
signal load_and_iterate_iterate_reg_1_cry_6 : std_logic;
signal \iterate_regZ0Z_0\ : std_logic;
signal iterate_reg_i_0 : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \iterate_regZ0Z_1\ : std_logic;
signal iterate_reg_i_1 : std_logic;
signal is_higher_than_un1_iterate_reg_cry_0 : std_logic;
signal \iterate_regZ0Z_2\ : std_logic;
signal iterate_reg_i_2 : std_logic;
signal is_higher_than_un1_iterate_reg_cry_1 : std_logic;
signal \iterate_regZ0Z_3\ : std_logic;
signal iterate_reg_i_3 : std_logic;
signal is_higher_than_un1_iterate_reg_cry_2 : std_logic;
signal \iterate_regZ0Z_4\ : std_logic;
signal iterate_reg_i_4 : std_logic;
signal is_higher_than_un1_iterate_reg_cry_3 : std_logic;
signal \iterate_regZ0Z_5\ : std_logic;
signal iterate_reg_i_5 : std_logic;
signal is_higher_than_un1_iterate_reg_cry_4 : std_logic;
signal \iterate_regZ0Z_6\ : std_logic;
signal iterate_reg_i_6 : std_logic;
signal is_higher_than_un1_iterate_reg_cry_5 : std_logic;
signal iterate_reg_i_7 : std_logic;
signal is_higher_than_un1_iterate_reg_cry_6 : std_logic;
signal iterate_ena_li : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \iterate_ena_li_THRU_CO_cascade_\ : std_logic;
signal \den_regZ0Z_5\ : std_logic;
signal \den_regZ0Z_6\ : std_logic;
signal \iterate_ena_li_THRU_CO\ : std_logic;
signal \counter_cntZ0Z_0\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \counter_cntZ0Z_1\ : std_logic;
signal counter_cnt_cry_0 : std_logic;
signal \counter_cntZ0Z_2\ : std_logic;
signal counter_cnt_cry_1 : std_logic;
signal \counter_cntZ0Z_3\ : std_logic;
signal counter_cnt_cry_2 : std_logic;
signal \counter_cntZ0Z_4\ : std_logic;
signal counter_cnt_cry_3 : std_logic;
signal \counter_cntZ0Z_5\ : std_logic;
signal counter_cnt_cry_4 : std_logic;
signal \counter_cntZ0Z_6\ : std_logic;
signal counter_cnt_cry_5 : std_logic;
signal counter_cnt_cry_6 : std_logic;
signal \counter_cntZ0Z_7\ : std_logic;
signal counter_cnte_0_i : std_logic;
signal \iterate_regZ0Z_7\ : std_logic;
signal load_and_iterate_iterate_reg_1_axb_7 : std_logic;
signal den_reg_i_3 : std_logic;
signal den_reg_i_4 : std_logic;
signal den_reg_i_1 : std_logic;
signal den_reg_i_2 : std_logic;
signal den_in_c_7 : std_logic;
signal \den_regZ0Z_7\ : std_logic;
signal den_in_c_2 : std_logic;
signal den_in_c_1 : std_logic;
signal den_in_c_3 : std_logic;
signal den_in_c_4 : std_logic;
signal \den_regZ0Z_4\ : std_logic;
signal \N_4_i\ : std_logic;
signal \den_regZ0Z_1\ : std_logic;
signal o2 : std_logic;
signal \den_regZ0Z_0\ : std_logic;
signal current_state_ns_i_sn_2 : std_logic;
signal is_den_zero_un5_den_reg_4 : std_logic;
signal current_state_ns_i_rn_1_2 : std_logic;
signal is_den_zero_un5_den_reg_3 : std_logic;
signal \resultOk_out_c\ : std_logic;
signal \divZero_out_c\ : std_logic;
signal \den_regZ0Z_3\ : std_logic;
signal \den_regZ0Z_2\ : std_logic;
signal m4_e_2 : std_logic;
signal \N_58_i\ : std_logic;
signal current_state_ns_i_0_1_0 : std_logic;
signal \current_stateZ0Z_5\ : std_logic;
signal \current_stateZ0Z_3\ : std_logic;
signal \N_60_2_c\ : std_logic;
signal \current_stateZ0Z_1\ : std_logic;
signal \current_stateZ0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_in_c_g : std_logic;
signal rst_in_n_c_i_g : std_logic;

signal clk_in_wire : std_logic;
signal den_in_wire : std_logic_vector(7 downto 0);
signal \divZero_out_wire\ : std_logic;
signal num_in_wire : std_logic_vector(7 downto 0);
signal res_out_wire : std_logic_vector(7 downto 0);
signal \resultOk_out_wire\ : std_logic;
signal rmn_out_wire : std_logic_vector(7 downto 0);
signal rst_in_n_wire : std_logic;
signal running_out_wire : std_logic;
signal start_in_wire : std_logic;

begin
    clk_in_wire <= clk_in;
    den_in_wire <= den_in;
    divZero_out <= \divZero_out_wire\;
    num_in_wire <= num_in;
    res_out <= res_out_wire;
    resultOk_out <= \resultOk_out_wire\;
    rmn_out <= rmn_out_wire;
    rst_in_n_wire <= rst_in_n;
    running_out <= running_out_wire;
    start_in_wire <= start_in;

    \clk_in_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__3512\,
            GLOBALBUFFEROUTPUT => clk_in_c_g
        );

    \clk_in_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3514\,
            DIN => \N__3513\,
            DOUT => \N__3512\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3514\,
            PADOUT => \N__3513\,
            PADIN => \N__3512\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \den_in_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3503\,
            DIN => \N__3502\,
            DOUT => \N__3501\,
            PACKAGEPIN => den_in_wire(0)
        );

    \den_in_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3503\,
            PADOUT => \N__3502\,
            PADIN => \N__3501\,
            CLOCKENABLE => 'H',
            DIN0 => den_in_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \den_in_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3494\,
            DIN => \N__3493\,
            DOUT => \N__3492\,
            PACKAGEPIN => den_in_wire(1)
        );

    \den_in_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3494\,
            PADOUT => \N__3493\,
            PADIN => \N__3492\,
            CLOCKENABLE => 'H',
            DIN0 => den_in_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \den_in_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3485\,
            DIN => \N__3484\,
            DOUT => \N__3483\,
            PACKAGEPIN => den_in_wire(2)
        );

    \den_in_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3485\,
            PADOUT => \N__3484\,
            PADIN => \N__3483\,
            CLOCKENABLE => 'H',
            DIN0 => den_in_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \den_in_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3476\,
            DIN => \N__3475\,
            DOUT => \N__3474\,
            PACKAGEPIN => den_in_wire(3)
        );

    \den_in_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3476\,
            PADOUT => \N__3475\,
            PADIN => \N__3474\,
            CLOCKENABLE => 'H',
            DIN0 => den_in_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \den_in_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3467\,
            DIN => \N__3466\,
            DOUT => \N__3465\,
            PACKAGEPIN => den_in_wire(4)
        );

    \den_in_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3467\,
            PADOUT => \N__3466\,
            PADIN => \N__3465\,
            CLOCKENABLE => 'H',
            DIN0 => den_in_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \den_in_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3458\,
            DIN => \N__3457\,
            DOUT => \N__3456\,
            PACKAGEPIN => den_in_wire(5)
        );

    \den_in_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3458\,
            PADOUT => \N__3457\,
            PADIN => \N__3456\,
            CLOCKENABLE => 'H',
            DIN0 => den_in_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \den_in_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3449\,
            DIN => \N__3448\,
            DOUT => \N__3447\,
            PACKAGEPIN => den_in_wire(6)
        );

    \den_in_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3449\,
            PADOUT => \N__3448\,
            PADIN => \N__3447\,
            CLOCKENABLE => 'H',
            DIN0 => den_in_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \den_in_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3440\,
            DIN => \N__3439\,
            DOUT => \N__3438\,
            PACKAGEPIN => den_in_wire(7)
        );

    \den_in_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3440\,
            PADOUT => \N__3439\,
            PADIN => \N__3438\,
            CLOCKENABLE => 'H',
            DIN0 => den_in_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \divZero_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3431\,
            DIN => \N__3430\,
            DOUT => \N__3429\,
            PACKAGEPIN => \divZero_out_wire\
        );

    \divZero_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3431\,
            PADOUT => \N__3430\,
            PADIN => \N__3429\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3133\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \num_in_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3422\,
            DIN => \N__3421\,
            DOUT => \N__3420\,
            PACKAGEPIN => num_in_wire(0)
        );

    \num_in_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3422\,
            PADOUT => \N__3421\,
            PADIN => \N__3420\,
            CLOCKENABLE => 'H',
            DIN0 => num_in_c_0,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \num_in_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3413\,
            DIN => \N__3412\,
            DOUT => \N__3411\,
            PACKAGEPIN => num_in_wire(1)
        );

    \num_in_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3413\,
            PADOUT => \N__3412\,
            PADIN => \N__3411\,
            CLOCKENABLE => 'H',
            DIN0 => num_in_c_1,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \num_in_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3404\,
            DIN => \N__3403\,
            DOUT => \N__3402\,
            PACKAGEPIN => num_in_wire(2)
        );

    \num_in_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3404\,
            PADOUT => \N__3403\,
            PADIN => \N__3402\,
            CLOCKENABLE => 'H',
            DIN0 => num_in_c_2,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \num_in_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3395\,
            DIN => \N__3394\,
            DOUT => \N__3393\,
            PACKAGEPIN => num_in_wire(3)
        );

    \num_in_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3395\,
            PADOUT => \N__3394\,
            PADIN => \N__3393\,
            CLOCKENABLE => 'H',
            DIN0 => num_in_c_3,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \num_in_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3386\,
            DIN => \N__3385\,
            DOUT => \N__3384\,
            PACKAGEPIN => num_in_wire(4)
        );

    \num_in_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3386\,
            PADOUT => \N__3385\,
            PADIN => \N__3384\,
            CLOCKENABLE => 'H',
            DIN0 => num_in_c_4,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \num_in_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3377\,
            DIN => \N__3376\,
            DOUT => \N__3375\,
            PACKAGEPIN => num_in_wire(5)
        );

    \num_in_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3377\,
            PADOUT => \N__3376\,
            PADIN => \N__3375\,
            CLOCKENABLE => 'H',
            DIN0 => num_in_c_5,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \num_in_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3368\,
            DIN => \N__3367\,
            DOUT => \N__3366\,
            PACKAGEPIN => num_in_wire(6)
        );

    \num_in_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3368\,
            PADOUT => \N__3367\,
            PADIN => \N__3366\,
            CLOCKENABLE => 'H',
            DIN0 => num_in_c_6,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \num_in_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3359\,
            DIN => \N__3358\,
            DOUT => \N__3357\,
            PACKAGEPIN => num_in_wire(7)
        );

    \num_in_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3359\,
            PADOUT => \N__3358\,
            PADIN => \N__3357\,
            CLOCKENABLE => 'H',
            DIN0 => num_in_c_7,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \res_out_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3350\,
            DIN => \N__3349\,
            DOUT => \N__3348\,
            PACKAGEPIN => res_out_wire(0)
        );

    \res_out_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3350\,
            PADOUT => \N__3349\,
            PADIN => \N__3348\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1747\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \res_out_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3341\,
            DIN => \N__3340\,
            DOUT => \N__3339\,
            PACKAGEPIN => res_out_wire(1)
        );

    \res_out_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3341\,
            PADOUT => \N__3340\,
            PADIN => \N__3339\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1861\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \res_out_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3332\,
            DIN => \N__3331\,
            DOUT => \N__3330\,
            PACKAGEPIN => res_out_wire(2)
        );

    \res_out_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3332\,
            PADOUT => \N__3331\,
            PADIN => \N__3330\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1891\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \res_out_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3323\,
            DIN => \N__3322\,
            DOUT => \N__3321\,
            PACKAGEPIN => res_out_wire(3)
        );

    \res_out_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3323\,
            PADOUT => \N__3322\,
            PADIN => \N__3321\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1726\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \res_out_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3314\,
            DIN => \N__3313\,
            DOUT => \N__3312\,
            PACKAGEPIN => res_out_wire(4)
        );

    \res_out_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3314\,
            PADOUT => \N__3313\,
            PADIN => \N__3312\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1909\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \res_out_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3305\,
            DIN => \N__3304\,
            DOUT => \N__3303\,
            PACKAGEPIN => res_out_wire(5)
        );

    \res_out_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3305\,
            PADOUT => \N__3304\,
            PADIN => \N__3303\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1873\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \res_out_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3296\,
            DIN => \N__3295\,
            DOUT => \N__3294\,
            PACKAGEPIN => res_out_wire(6)
        );

    \res_out_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3296\,
            PADOUT => \N__3295\,
            PADIN => \N__3294\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1693\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \res_out_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3287\,
            DIN => \N__3286\,
            DOUT => \N__3285\,
            PACKAGEPIN => res_out_wire(7)
        );

    \res_out_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3287\,
            PADOUT => \N__3286\,
            PADIN => \N__3285\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1708\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \resultOk_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3278\,
            DIN => \N__3277\,
            DOUT => \N__3276\,
            PACKAGEPIN => \resultOk_out_wire\
        );

    \resultOk_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3278\,
            PADOUT => \N__3277\,
            PADIN => \N__3276\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3160\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rmn_out_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3269\,
            DIN => \N__3268\,
            DOUT => \N__3267\,
            PACKAGEPIN => rmn_out_wire(0)
        );

    \rmn_out_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3269\,
            PADOUT => \N__3268\,
            PADIN => \N__3267\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1786\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rmn_out_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3260\,
            DIN => \N__3259\,
            DOUT => \N__3258\,
            PACKAGEPIN => rmn_out_wire(1)
        );

    \rmn_out_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3260\,
            PADOUT => \N__3259\,
            PADIN => \N__3258\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1762\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rmn_out_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3251\,
            DIN => \N__3250\,
            DOUT => \N__3249\,
            PACKAGEPIN => rmn_out_wire(2)
        );

    \rmn_out_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3251\,
            PADOUT => \N__3250\,
            PADIN => \N__3249\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1771\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rmn_out_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3242\,
            DIN => \N__3241\,
            DOUT => \N__3240\,
            PACKAGEPIN => rmn_out_wire(3)
        );

    \rmn_out_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3242\,
            PADOUT => \N__3241\,
            PADIN => \N__3240\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1567\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rmn_out_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3233\,
            DIN => \N__3232\,
            DOUT => \N__3231\,
            PACKAGEPIN => rmn_out_wire(4)
        );

    \rmn_out_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3233\,
            PADOUT => \N__3232\,
            PADIN => \N__3231\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1558\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rmn_out_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3224\,
            DIN => \N__3223\,
            DOUT => \N__3222\,
            PACKAGEPIN => rmn_out_wire(5)
        );

    \rmn_out_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3224\,
            PADOUT => \N__3223\,
            PADIN => \N__3222\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1816\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rmn_out_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3215\,
            DIN => \N__3214\,
            DOUT => \N__3213\,
            PACKAGEPIN => rmn_out_wire(6)
        );

    \rmn_out_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3215\,
            PADOUT => \N__3214\,
            PADIN => \N__3213\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1801\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rmn_out_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3206\,
            DIN => \N__3205\,
            DOUT => \N__3204\,
            PACKAGEPIN => rmn_out_wire(7)
        );

    \rmn_out_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3206\,
            PADOUT => \N__3205\,
            PADIN => \N__3204\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__1585\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \rst_in_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3197\,
            DIN => \N__3196\,
            DOUT => \N__3195\,
            PACKAGEPIN => rst_in_n_wire
        );

    \rst_in_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3197\,
            PADOUT => \N__3196\,
            PADIN => \N__3195\,
            CLOCKENABLE => 'H',
            DIN0 => rst_in_n_c,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \running_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3188\,
            DIN => \N__3187\,
            DOUT => \N__3186\,
            PACKAGEPIN => running_out_wire
        );

    \running_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__3188\,
            PADOUT => \N__3187\,
            PADIN => \N__3186\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__3043\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \start_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__3179\,
            DIN => \N__3178\,
            DOUT => \N__3177\,
            PACKAGEPIN => start_in_wire
        );

    \start_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__3179\,
            PADOUT => \N__3178\,
            PADIN => \N__3177\,
            CLOCKENABLE => 'H',
            DIN0 => \N_60_2_c\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__698\ : IoInMux
    port map (
            O => \N__3160\,
            I => \N__3157\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3157\,
            I => \N__3154\
        );

    \I__696\ : Span4Mux_s2_h
    port map (
            O => \N__3154\,
            I => \N__3151\
        );

    \I__695\ : Span4Mux_v
    port map (
            O => \N__3151\,
            I => \N__3147\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__3150\,
            I => \N__3144\
        );

    \I__693\ : Span4Mux_h
    port map (
            O => \N__3147\,
            I => \N__3141\
        );

    \I__692\ : InMux
    port map (
            O => \N__3144\,
            I => \N__3138\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__3141\,
            I => \resultOk_out_c\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__3138\,
            I => \resultOk_out_c\
        );

    \I__689\ : IoInMux
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3130\,
            I => \N__3127\
        );

    \I__687\ : IoSpan4Mux
    port map (
            O => \N__3127\,
            I => \N__3124\
        );

    \I__686\ : IoSpan4Mux
    port map (
            O => \N__3124\,
            I => \N__3121\
        );

    \I__685\ : Span4Mux_s3_h
    port map (
            O => \N__3121\,
            I => \N__3117\
        );

    \I__684\ : InMux
    port map (
            O => \N__3120\,
            I => \N__3114\
        );

    \I__683\ : Odrv4
    port map (
            O => \N__3117\,
            I => \divZero_out_c\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3114\,
            I => \divZero_out_c\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__3109\,
            I => \N__3104\
        );

    \I__680\ : InMux
    port map (
            O => \N__3108\,
            I => \N__3101\
        );

    \I__679\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3097\
        );

    \I__678\ : InMux
    port map (
            O => \N__3104\,
            I => \N__3094\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3101\,
            I => \N__3091\
        );

    \I__676\ : InMux
    port map (
            O => \N__3100\,
            I => \N__3088\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3097\,
            I => \N__3085\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3094\,
            I => \den_regZ0Z_3\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__3091\,
            I => \den_regZ0Z_3\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3088\,
            I => \den_regZ0Z_3\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__3085\,
            I => \den_regZ0Z_3\
        );

    \I__670\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3072\
        );

    \I__669\ : InMux
    port map (
            O => \N__3075\,
            I => \N__3067\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3072\,
            I => \N__3064\
        );

    \I__667\ : InMux
    port map (
            O => \N__3071\,
            I => \N__3061\
        );

    \I__666\ : InMux
    port map (
            O => \N__3070\,
            I => \N__3058\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3067\,
            I => \den_regZ0Z_2\
        );

    \I__664\ : Odrv4
    port map (
            O => \N__3064\,
            I => \den_regZ0Z_2\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3061\,
            I => \den_regZ0Z_2\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3058\,
            I => \den_regZ0Z_2\
        );

    \I__661\ : InMux
    port map (
            O => \N__3049\,
            I => \N__3046\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3046\,
            I => m4_e_2
        );

    \I__659\ : IoInMux
    port map (
            O => \N__3043\,
            I => \N__3040\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3040\,
            I => \N__3037\
        );

    \I__657\ : Span4Mux_s3_h
    port map (
            O => \N__3037\,
            I => \N__3034\
        );

    \I__656\ : Span4Mux_v
    port map (
            O => \N__3034\,
            I => \N__3031\
        );

    \I__655\ : Span4Mux_v
    port map (
            O => \N__3031\,
            I => \N__3028\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__3028\,
            I => \N_58_i\
        );

    \I__653\ : InMux
    port map (
            O => \N__3025\,
            I => \N__3022\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3022\,
            I => \N__3019\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__3019\,
            I => current_state_ns_i_0_1_0
        );

    \I__650\ : InMux
    port map (
            O => \N__3016\,
            I => \N__3012\
        );

    \I__649\ : InMux
    port map (
            O => \N__3015\,
            I => \N__3009\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3012\,
            I => \current_stateZ0Z_5\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3009\,
            I => \current_stateZ0Z_5\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__3004\,
            I => \N__3000\
        );

    \I__645\ : InMux
    port map (
            O => \N__3003\,
            I => \N__2995\
        );

    \I__644\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2990\
        );

    \I__643\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2990\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__2998\,
            I => \N__2986\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__2995\,
            I => \N__2979\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__2990\,
            I => \N__2979\
        );

    \I__639\ : InMux
    port map (
            O => \N__2989\,
            I => \N__2974\
        );

    \I__638\ : InMux
    port map (
            O => \N__2986\,
            I => \N__2974\
        );

    \I__637\ : InMux
    port map (
            O => \N__2985\,
            I => \N__2969\
        );

    \I__636\ : InMux
    port map (
            O => \N__2984\,
            I => \N__2969\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__2979\,
            I => \current_stateZ0Z_3\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__2974\,
            I => \current_stateZ0Z_3\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__2969\,
            I => \current_stateZ0Z_3\
        );

    \I__632\ : InMux
    port map (
            O => \N__2962\,
            I => \N__2958\
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__2961\,
            I => \N__2954\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__2958\,
            I => \N__2951\
        );

    \I__629\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2946\
        );

    \I__628\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2946\
        );

    \I__627\ : Span4Mux_h
    port map (
            O => \N__2951\,
            I => \N__2941\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__2946\,
            I => \N__2941\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__2941\,
            I => \N__2938\
        );

    \I__624\ : Sp12to4
    port map (
            O => \N__2938\,
            I => \N__2935\
        );

    \I__623\ : Odrv12
    port map (
            O => \N__2935\,
            I => \N_60_2_c\
        );

    \I__622\ : InMux
    port map (
            O => \N__2932\,
            I => \N__2926\
        );

    \I__621\ : InMux
    port map (
            O => \N__2931\,
            I => \N__2926\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__2926\,
            I => \N__2919\
        );

    \I__619\ : InMux
    port map (
            O => \N__2925\,
            I => \N__2914\
        );

    \I__618\ : InMux
    port map (
            O => \N__2924\,
            I => \N__2914\
        );

    \I__617\ : InMux
    port map (
            O => \N__2923\,
            I => \N__2911\
        );

    \I__616\ : InMux
    port map (
            O => \N__2922\,
            I => \N__2908\
        );

    \I__615\ : Odrv4
    port map (
            O => \N__2919\,
            I => \current_stateZ0Z_1\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__2914\,
            I => \current_stateZ0Z_1\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__2911\,
            I => \current_stateZ0Z_1\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__2908\,
            I => \current_stateZ0Z_1\
        );

    \I__611\ : CEMux
    port map (
            O => \N__2899\,
            I => \N__2887\
        );

    \I__610\ : InMux
    port map (
            O => \N__2898\,
            I => \N__2872\
        );

    \I__609\ : InMux
    port map (
            O => \N__2897\,
            I => \N__2872\
        );

    \I__608\ : InMux
    port map (
            O => \N__2896\,
            I => \N__2872\
        );

    \I__607\ : InMux
    port map (
            O => \N__2895\,
            I => \N__2872\
        );

    \I__606\ : InMux
    port map (
            O => \N__2894\,
            I => \N__2872\
        );

    \I__605\ : InMux
    port map (
            O => \N__2893\,
            I => \N__2872\
        );

    \I__604\ : InMux
    port map (
            O => \N__2892\,
            I => \N__2872\
        );

    \I__603\ : CEMux
    port map (
            O => \N__2891\,
            I => \N__2868\
        );

    \I__602\ : InMux
    port map (
            O => \N__2890\,
            I => \N__2865\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__2887\,
            I => \N__2853\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__2872\,
            I => \N__2850\
        );

    \I__599\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2847\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__2868\,
            I => \N__2842\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__2865\,
            I => \N__2842\
        );

    \I__596\ : InMux
    port map (
            O => \N__2864\,
            I => \N__2839\
        );

    \I__595\ : InMux
    port map (
            O => \N__2863\,
            I => \N__2828\
        );

    \I__594\ : InMux
    port map (
            O => \N__2862\,
            I => \N__2828\
        );

    \I__593\ : InMux
    port map (
            O => \N__2861\,
            I => \N__2828\
        );

    \I__592\ : InMux
    port map (
            O => \N__2860\,
            I => \N__2828\
        );

    \I__591\ : InMux
    port map (
            O => \N__2859\,
            I => \N__2828\
        );

    \I__590\ : InMux
    port map (
            O => \N__2858\,
            I => \N__2821\
        );

    \I__589\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2821\
        );

    \I__588\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2821\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__2853\,
            I => \N__2818\
        );

    \I__586\ : Span4Mux_v
    port map (
            O => \N__2850\,
            I => \N__2815\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__2847\,
            I => \N__2808\
        );

    \I__584\ : Span4Mux_h
    port map (
            O => \N__2842\,
            I => \N__2808\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__2839\,
            I => \N__2808\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__2828\,
            I => \current_stateZ0Z_0\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__2821\,
            I => \current_stateZ0Z_0\
        );

    \I__580\ : Odrv4
    port map (
            O => \N__2818\,
            I => \current_stateZ0Z_0\
        );

    \I__579\ : Odrv4
    port map (
            O => \N__2815\,
            I => \current_stateZ0Z_0\
        );

    \I__578\ : Odrv4
    port map (
            O => \N__2808\,
            I => \current_stateZ0Z_0\
        );

    \I__577\ : ClkMux
    port map (
            O => \N__2797\,
            I => \N__2770\
        );

    \I__576\ : ClkMux
    port map (
            O => \N__2796\,
            I => \N__2770\
        );

    \I__575\ : ClkMux
    port map (
            O => \N__2795\,
            I => \N__2770\
        );

    \I__574\ : ClkMux
    port map (
            O => \N__2794\,
            I => \N__2770\
        );

    \I__573\ : ClkMux
    port map (
            O => \N__2793\,
            I => \N__2770\
        );

    \I__572\ : ClkMux
    port map (
            O => \N__2792\,
            I => \N__2770\
        );

    \I__571\ : ClkMux
    port map (
            O => \N__2791\,
            I => \N__2770\
        );

    \I__570\ : ClkMux
    port map (
            O => \N__2790\,
            I => \N__2770\
        );

    \I__569\ : ClkMux
    port map (
            O => \N__2789\,
            I => \N__2770\
        );

    \I__568\ : GlobalMux
    port map (
            O => \N__2770\,
            I => \N__2767\
        );

    \I__567\ : gio2CtrlBuf
    port map (
            O => \N__2767\,
            I => clk_in_c_g
        );

    \I__566\ : SRMux
    port map (
            O => \N__2764\,
            I => \N__2737\
        );

    \I__565\ : SRMux
    port map (
            O => \N__2763\,
            I => \N__2737\
        );

    \I__564\ : SRMux
    port map (
            O => \N__2762\,
            I => \N__2737\
        );

    \I__563\ : SRMux
    port map (
            O => \N__2761\,
            I => \N__2737\
        );

    \I__562\ : SRMux
    port map (
            O => \N__2760\,
            I => \N__2737\
        );

    \I__561\ : SRMux
    port map (
            O => \N__2759\,
            I => \N__2737\
        );

    \I__560\ : SRMux
    port map (
            O => \N__2758\,
            I => \N__2737\
        );

    \I__559\ : SRMux
    port map (
            O => \N__2757\,
            I => \N__2737\
        );

    \I__558\ : SRMux
    port map (
            O => \N__2756\,
            I => \N__2737\
        );

    \I__557\ : GlobalMux
    port map (
            O => \N__2737\,
            I => \N__2734\
        );

    \I__556\ : gio2CtrlBuf
    port map (
            O => \N__2734\,
            I => rst_in_n_c_i_g
        );

    \I__555\ : InMux
    port map (
            O => \N__2731\,
            I => \N__2728\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__2728\,
            I => \N__2725\
        );

    \I__553\ : Span4Mux_v
    port map (
            O => \N__2725\,
            I => \N__2722\
        );

    \I__552\ : Sp12to4
    port map (
            O => \N__2722\,
            I => \N__2719\
        );

    \I__551\ : Span12Mux_h
    port map (
            O => \N__2719\,
            I => \N__2716\
        );

    \I__550\ : Span12Mux_v
    port map (
            O => \N__2716\,
            I => \N__2713\
        );

    \I__549\ : Odrv12
    port map (
            O => \N__2713\,
            I => den_in_c_2
        );

    \I__548\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2707\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__2707\,
            I => \N__2704\
        );

    \I__546\ : Span4Mux_v
    port map (
            O => \N__2704\,
            I => \N__2701\
        );

    \I__545\ : Span4Mux_h
    port map (
            O => \N__2701\,
            I => \N__2698\
        );

    \I__544\ : Sp12to4
    port map (
            O => \N__2698\,
            I => \N__2695\
        );

    \I__543\ : Span12Mux_v
    port map (
            O => \N__2695\,
            I => \N__2692\
        );

    \I__542\ : Odrv12
    port map (
            O => \N__2692\,
            I => den_in_c_1
        );

    \I__541\ : InMux
    port map (
            O => \N__2689\,
            I => \N__2686\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2686\,
            I => \N__2683\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__2683\,
            I => \N__2680\
        );

    \I__538\ : Span4Mux_h
    port map (
            O => \N__2680\,
            I => \N__2677\
        );

    \I__537\ : Span4Mux_v
    port map (
            O => \N__2677\,
            I => \N__2674\
        );

    \I__536\ : Span4Mux_v
    port map (
            O => \N__2674\,
            I => \N__2671\
        );

    \I__535\ : Odrv4
    port map (
            O => \N__2671\,
            I => den_in_c_3
        );

    \I__534\ : InMux
    port map (
            O => \N__2668\,
            I => \N__2665\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__2665\,
            I => \N__2662\
        );

    \I__532\ : Sp12to4
    port map (
            O => \N__2662\,
            I => \N__2659\
        );

    \I__531\ : Span12Mux_v
    port map (
            O => \N__2659\,
            I => \N__2656\
        );

    \I__530\ : Odrv12
    port map (
            O => \N__2656\,
            I => den_in_c_4
        );

    \I__529\ : InMux
    port map (
            O => \N__2653\,
            I => \N__2645\
        );

    \I__528\ : InMux
    port map (
            O => \N__2652\,
            I => \N__2645\
        );

    \I__527\ : InMux
    port map (
            O => \N__2651\,
            I => \N__2642\
        );

    \I__526\ : InMux
    port map (
            O => \N__2650\,
            I => \N__2639\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__2645\,
            I => \den_regZ0Z_4\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__2642\,
            I => \den_regZ0Z_4\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__2639\,
            I => \den_regZ0Z_4\
        );

    \I__522\ : CEMux
    port map (
            O => \N__2632\,
            I => \N__2627\
        );

    \I__521\ : CEMux
    port map (
            O => \N__2631\,
            I => \N__2624\
        );

    \I__520\ : InMux
    port map (
            O => \N__2630\,
            I => \N__2621\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__2627\,
            I => \N_4_i\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__2624\,
            I => \N_4_i\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__2621\,
            I => \N_4_i\
        );

    \I__516\ : InMux
    port map (
            O => \N__2614\,
            I => \N__2608\
        );

    \I__515\ : InMux
    port map (
            O => \N__2613\,
            I => \N__2605\
        );

    \I__514\ : InMux
    port map (
            O => \N__2612\,
            I => \N__2602\
        );

    \I__513\ : InMux
    port map (
            O => \N__2611\,
            I => \N__2599\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__2608\,
            I => \den_regZ0Z_1\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__2605\,
            I => \den_regZ0Z_1\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__2602\,
            I => \den_regZ0Z_1\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__2599\,
            I => \den_regZ0Z_1\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__2590\,
            I => \N__2587\
        );

    \I__507\ : InMux
    port map (
            O => \N__2587\,
            I => \N__2584\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__2584\,
            I => o2
        );

    \I__505\ : InMux
    port map (
            O => \N__2581\,
            I => \N__2578\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__2578\,
            I => \N__2573\
        );

    \I__503\ : InMux
    port map (
            O => \N__2577\,
            I => \N__2570\
        );

    \I__502\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2565\
        );

    \I__501\ : Span4Mux_h
    port map (
            O => \N__2573\,
            I => \N__2560\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2570\,
            I => \N__2560\
        );

    \I__499\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2557\
        );

    \I__498\ : InMux
    port map (
            O => \N__2568\,
            I => \N__2554\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__2565\,
            I => \den_regZ0Z_0\
        );

    \I__496\ : Odrv4
    port map (
            O => \N__2560\,
            I => \den_regZ0Z_0\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__2557\,
            I => \den_regZ0Z_0\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__2554\,
            I => \den_regZ0Z_0\
        );

    \I__493\ : InMux
    port map (
            O => \N__2545\,
            I => \N__2542\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__2542\,
            I => current_state_ns_i_sn_2
        );

    \I__491\ : InMux
    port map (
            O => \N__2539\,
            I => \N__2536\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2536\,
            I => is_den_zero_un5_den_reg_4
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__2533\,
            I => \N__2530\
        );

    \I__488\ : InMux
    port map (
            O => \N__2530\,
            I => \N__2527\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__2527\,
            I => current_state_ns_i_rn_1_2
        );

    \I__486\ : InMux
    port map (
            O => \N__2524\,
            I => \N__2521\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__2521\,
            I => is_den_zero_un5_den_reg_3
        );

    \I__484\ : InMux
    port map (
            O => \N__2518\,
            I => \N__2514\
        );

    \I__483\ : InMux
    port map (
            O => \N__2517\,
            I => \N__2511\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__2514\,
            I => \counter_cntZ0Z_5\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2511\,
            I => \counter_cntZ0Z_5\
        );

    \I__480\ : InMux
    port map (
            O => \N__2506\,
            I => counter_cnt_cry_4
        );

    \I__479\ : InMux
    port map (
            O => \N__2503\,
            I => \N__2499\
        );

    \I__478\ : InMux
    port map (
            O => \N__2502\,
            I => \N__2496\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__2499\,
            I => \counter_cntZ0Z_6\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2496\,
            I => \counter_cntZ0Z_6\
        );

    \I__475\ : InMux
    port map (
            O => \N__2491\,
            I => counter_cnt_cry_5
        );

    \I__474\ : InMux
    port map (
            O => \N__2488\,
            I => counter_cnt_cry_6
        );

    \I__473\ : InMux
    port map (
            O => \N__2485\,
            I => \N__2481\
        );

    \I__472\ : InMux
    port map (
            O => \N__2484\,
            I => \N__2478\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__2481\,
            I => \counter_cntZ0Z_7\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__2478\,
            I => \counter_cntZ0Z_7\
        );

    \I__469\ : CEMux
    port map (
            O => \N__2473\,
            I => \N__2469\
        );

    \I__468\ : CEMux
    port map (
            O => \N__2472\,
            I => \N__2465\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__2469\,
            I => \N__2462\
        );

    \I__466\ : CEMux
    port map (
            O => \N__2468\,
            I => \N__2459\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__2465\,
            I => \N__2456\
        );

    \I__464\ : Span4Mux_v
    port map (
            O => \N__2462\,
            I => \N__2451\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2459\,
            I => \N__2451\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__2456\,
            I => counter_cnte_0_i
        );

    \I__461\ : Odrv4
    port map (
            O => \N__2451\,
            I => counter_cnte_0_i
        );

    \I__460\ : InMux
    port map (
            O => \N__2446\,
            I => \N__2443\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2443\,
            I => \N__2438\
        );

    \I__458\ : InMux
    port map (
            O => \N__2442\,
            I => \N__2435\
        );

    \I__457\ : InMux
    port map (
            O => \N__2441\,
            I => \N__2432\
        );

    \I__456\ : Odrv4
    port map (
            O => \N__2438\,
            I => \iterate_regZ0Z_7\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2435\,
            I => \iterate_regZ0Z_7\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__2432\,
            I => \iterate_regZ0Z_7\
        );

    \I__453\ : InMux
    port map (
            O => \N__2425\,
            I => \N__2422\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2422\,
            I => load_and_iterate_iterate_reg_1_axb_7
        );

    \I__451\ : CascadeMux
    port map (
            O => \N__2419\,
            I => \N__2416\
        );

    \I__450\ : InMux
    port map (
            O => \N__2416\,
            I => \N__2413\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2413\,
            I => den_reg_i_3
        );

    \I__448\ : InMux
    port map (
            O => \N__2410\,
            I => \N__2407\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2407\,
            I => den_reg_i_4
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__2404\,
            I => \N__2401\
        );

    \I__445\ : InMux
    port map (
            O => \N__2401\,
            I => \N__2398\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2398\,
            I => den_reg_i_1
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__2395\,
            I => \N__2392\
        );

    \I__442\ : InMux
    port map (
            O => \N__2392\,
            I => \N__2389\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2389\,
            I => den_reg_i_2
        );

    \I__440\ : InMux
    port map (
            O => \N__2386\,
            I => \N__2383\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2383\,
            I => \N__2380\
        );

    \I__438\ : Sp12to4
    port map (
            O => \N__2380\,
            I => \N__2377\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__2377\,
            I => \N__2374\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__2374\,
            I => den_in_c_7
        );

    \I__435\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2363\
        );

    \I__434\ : InMux
    port map (
            O => \N__2370\,
            I => \N__2363\
        );

    \I__433\ : InMux
    port map (
            O => \N__2369\,
            I => \N__2360\
        );

    \I__432\ : InMux
    port map (
            O => \N__2368\,
            I => \N__2357\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2363\,
            I => \den_regZ0Z_7\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2360\,
            I => \den_regZ0Z_7\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2357\,
            I => \den_regZ0Z_7\
        );

    \I__428\ : CascadeMux
    port map (
            O => \N__2350\,
            I => \N__2347\
        );

    \I__427\ : InMux
    port map (
            O => \N__2347\,
            I => \N__2339\
        );

    \I__426\ : InMux
    port map (
            O => \N__2346\,
            I => \N__2339\
        );

    \I__425\ : InMux
    port map (
            O => \N__2345\,
            I => \N__2336\
        );

    \I__424\ : InMux
    port map (
            O => \N__2344\,
            I => \N__2333\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2339\,
            I => \N__2328\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2336\,
            I => \N__2328\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2333\,
            I => \den_regZ0Z_5\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__2328\,
            I => \den_regZ0Z_5\
        );

    \I__419\ : InMux
    port map (
            O => \N__2323\,
            I => \N__2319\
        );

    \I__418\ : InMux
    port map (
            O => \N__2322\,
            I => \N__2316\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2319\,
            I => \N__2311\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__2316\,
            I => \N__2311\
        );

    \I__415\ : Span4Mux_h
    port map (
            O => \N__2311\,
            I => \N__2306\
        );

    \I__414\ : InMux
    port map (
            O => \N__2310\,
            I => \N__2303\
        );

    \I__413\ : InMux
    port map (
            O => \N__2309\,
            I => \N__2300\
        );

    \I__412\ : Odrv4
    port map (
            O => \N__2306\,
            I => \den_regZ0Z_6\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2303\,
            I => \den_regZ0Z_6\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2300\,
            I => \den_regZ0Z_6\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__2293\,
            I => \N__2290\
        );

    \I__408\ : InMux
    port map (
            O => \N__2290\,
            I => \N__2284\
        );

    \I__407\ : InMux
    port map (
            O => \N__2289\,
            I => \N__2284\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2284\,
            I => \iterate_ena_li_THRU_CO\
        );

    \I__405\ : InMux
    port map (
            O => \N__2281\,
            I => \N__2277\
        );

    \I__404\ : InMux
    port map (
            O => \N__2280\,
            I => \N__2274\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2277\,
            I => \counter_cntZ0Z_0\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2274\,
            I => \counter_cntZ0Z_0\
        );

    \I__401\ : InMux
    port map (
            O => \N__2269\,
            I => \bfn_2_13_0_\
        );

    \I__400\ : InMux
    port map (
            O => \N__2266\,
            I => \N__2262\
        );

    \I__399\ : InMux
    port map (
            O => \N__2265\,
            I => \N__2259\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2262\,
            I => \counter_cntZ0Z_1\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2259\,
            I => \counter_cntZ0Z_1\
        );

    \I__396\ : InMux
    port map (
            O => \N__2254\,
            I => counter_cnt_cry_0
        );

    \I__395\ : InMux
    port map (
            O => \N__2251\,
            I => \N__2247\
        );

    \I__394\ : InMux
    port map (
            O => \N__2250\,
            I => \N__2244\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2247\,
            I => \counter_cntZ0Z_2\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2244\,
            I => \counter_cntZ0Z_2\
        );

    \I__391\ : InMux
    port map (
            O => \N__2239\,
            I => counter_cnt_cry_1
        );

    \I__390\ : InMux
    port map (
            O => \N__2236\,
            I => \N__2232\
        );

    \I__389\ : InMux
    port map (
            O => \N__2235\,
            I => \N__2229\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2232\,
            I => \counter_cntZ0Z_3\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2229\,
            I => \counter_cntZ0Z_3\
        );

    \I__386\ : InMux
    port map (
            O => \N__2224\,
            I => counter_cnt_cry_2
        );

    \I__385\ : InMux
    port map (
            O => \N__2221\,
            I => \N__2217\
        );

    \I__384\ : InMux
    port map (
            O => \N__2220\,
            I => \N__2214\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2217\,
            I => \counter_cntZ0Z_4\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2214\,
            I => \counter_cntZ0Z_4\
        );

    \I__381\ : InMux
    port map (
            O => \N__2209\,
            I => counter_cnt_cry_3
        );

    \I__380\ : CascadeMux
    port map (
            O => \N__2206\,
            I => \N__2203\
        );

    \I__379\ : InMux
    port map (
            O => \N__2203\,
            I => \N__2200\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2200\,
            I => iterate_reg_i_3
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__2197\,
            I => \N__2193\
        );

    \I__376\ : InMux
    port map (
            O => \N__2196\,
            I => \N__2189\
        );

    \I__375\ : InMux
    port map (
            O => \N__2193\,
            I => \N__2186\
        );

    \I__374\ : InMux
    port map (
            O => \N__2192\,
            I => \N__2183\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2189\,
            I => \iterate_regZ0Z_4\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2186\,
            I => \iterate_regZ0Z_4\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2183\,
            I => \iterate_regZ0Z_4\
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__2176\,
            I => \N__2173\
        );

    \I__369\ : InMux
    port map (
            O => \N__2173\,
            I => \N__2170\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2170\,
            I => iterate_reg_i_4
        );

    \I__367\ : InMux
    port map (
            O => \N__2167\,
            I => \N__2162\
        );

    \I__366\ : InMux
    port map (
            O => \N__2166\,
            I => \N__2159\
        );

    \I__365\ : InMux
    port map (
            O => \N__2165\,
            I => \N__2156\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2162\,
            I => \iterate_regZ0Z_5\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2159\,
            I => \iterate_regZ0Z_5\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2156\,
            I => \iterate_regZ0Z_5\
        );

    \I__361\ : CascadeMux
    port map (
            O => \N__2149\,
            I => \N__2146\
        );

    \I__360\ : InMux
    port map (
            O => \N__2146\,
            I => \N__2143\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2143\,
            I => iterate_reg_i_5
        );

    \I__358\ : InMux
    port map (
            O => \N__2140\,
            I => \N__2135\
        );

    \I__357\ : InMux
    port map (
            O => \N__2139\,
            I => \N__2132\
        );

    \I__356\ : InMux
    port map (
            O => \N__2138\,
            I => \N__2129\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2135\,
            I => \iterate_regZ0Z_6\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2132\,
            I => \iterate_regZ0Z_6\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2129\,
            I => \iterate_regZ0Z_6\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__2122\,
            I => \N__2119\
        );

    \I__351\ : InMux
    port map (
            O => \N__2119\,
            I => \N__2116\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2116\,
            I => iterate_reg_i_6
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__2113\,
            I => \N__2110\
        );

    \I__348\ : InMux
    port map (
            O => \N__2110\,
            I => \N__2107\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2107\,
            I => iterate_reg_i_7
        );

    \I__346\ : InMux
    port map (
            O => \N__2104\,
            I => \bfn_2_12_0_\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__2101\,
            I => \iterate_ena_li_THRU_CO_cascade_\
        );

    \I__344\ : InMux
    port map (
            O => \N__2098\,
            I => \N__2095\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2095\,
            I => load_and_iterate_iterate_reg_1_3
        );

    \I__342\ : InMux
    port map (
            O => \N__2092\,
            I => load_and_iterate_iterate_reg_1_cry_2
        );

    \I__341\ : InMux
    port map (
            O => \N__2089\,
            I => \N__2086\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2086\,
            I => load_and_iterate_iterate_reg_1_4
        );

    \I__339\ : InMux
    port map (
            O => \N__2083\,
            I => load_and_iterate_iterate_reg_1_cry_3
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__2080\,
            I => \N__2077\
        );

    \I__337\ : InMux
    port map (
            O => \N__2077\,
            I => \N__2074\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2074\,
            I => den_reg_i_5
        );

    \I__335\ : InMux
    port map (
            O => \N__2071\,
            I => \N__2068\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2068\,
            I => load_and_iterate_iterate_reg_1_5
        );

    \I__333\ : InMux
    port map (
            O => \N__2065\,
            I => load_and_iterate_iterate_reg_1_cry_4
        );

    \I__332\ : CascadeMux
    port map (
            O => \N__2062\,
            I => \N__2059\
        );

    \I__331\ : InMux
    port map (
            O => \N__2059\,
            I => \N__2056\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2056\,
            I => den_reg_i_6
        );

    \I__329\ : InMux
    port map (
            O => \N__2053\,
            I => \N__2050\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2050\,
            I => load_and_iterate_iterate_reg_1_6
        );

    \I__327\ : InMux
    port map (
            O => \N__2047\,
            I => load_and_iterate_iterate_reg_1_cry_5
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__2044\,
            I => \N__2041\
        );

    \I__325\ : InMux
    port map (
            O => \N__2041\,
            I => \N__2038\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2038\,
            I => \N__2035\
        );

    \I__323\ : Span4Mux_v
    port map (
            O => \N__2035\,
            I => \N__2032\
        );

    \I__322\ : Span4Mux_v
    port map (
            O => \N__2032\,
            I => \N__2029\
        );

    \I__321\ : Span4Mux_v
    port map (
            O => \N__2029\,
            I => \N__2026\
        );

    \I__320\ : Span4Mux_v
    port map (
            O => \N__2026\,
            I => \N__2023\
        );

    \I__319\ : IoSpan4Mux
    port map (
            O => \N__2023\,
            I => \N__2020\
        );

    \I__318\ : Odrv4
    port map (
            O => \N__2020\,
            I => num_in_c_7
        );

    \I__317\ : InMux
    port map (
            O => \N__2017\,
            I => load_and_iterate_iterate_reg_1_cry_6
        );

    \I__316\ : InMux
    port map (
            O => \N__2014\,
            I => \N__2008\
        );

    \I__315\ : InMux
    port map (
            O => \N__2013\,
            I => \N__2005\
        );

    \I__314\ : InMux
    port map (
            O => \N__2012\,
            I => \N__2002\
        );

    \I__313\ : InMux
    port map (
            O => \N__2011\,
            I => \N__1999\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2008\,
            I => \iterate_regZ0Z_0\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2005\,
            I => \iterate_regZ0Z_0\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2002\,
            I => \iterate_regZ0Z_0\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__1999\,
            I => \iterate_regZ0Z_0\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__1990\,
            I => \N__1987\
        );

    \I__307\ : InMux
    port map (
            O => \N__1987\,
            I => \N__1984\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__1984\,
            I => iterate_reg_i_0
        );

    \I__305\ : InMux
    port map (
            O => \N__1981\,
            I => \N__1976\
        );

    \I__304\ : InMux
    port map (
            O => \N__1980\,
            I => \N__1973\
        );

    \I__303\ : InMux
    port map (
            O => \N__1979\,
            I => \N__1970\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__1976\,
            I => \iterate_regZ0Z_1\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__1973\,
            I => \iterate_regZ0Z_1\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1970\,
            I => \iterate_regZ0Z_1\
        );

    \I__299\ : CascadeMux
    port map (
            O => \N__1963\,
            I => \N__1960\
        );

    \I__298\ : InMux
    port map (
            O => \N__1960\,
            I => \N__1957\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__1957\,
            I => iterate_reg_i_1
        );

    \I__296\ : InMux
    port map (
            O => \N__1954\,
            I => \N__1949\
        );

    \I__295\ : InMux
    port map (
            O => \N__1953\,
            I => \N__1946\
        );

    \I__294\ : InMux
    port map (
            O => \N__1952\,
            I => \N__1943\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__1949\,
            I => \iterate_regZ0Z_2\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1946\,
            I => \iterate_regZ0Z_2\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__1943\,
            I => \iterate_regZ0Z_2\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__1936\,
            I => \N__1933\
        );

    \I__289\ : InMux
    port map (
            O => \N__1933\,
            I => \N__1930\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__1930\,
            I => iterate_reg_i_2
        );

    \I__287\ : InMux
    port map (
            O => \N__1927\,
            I => \N__1922\
        );

    \I__286\ : InMux
    port map (
            O => \N__1926\,
            I => \N__1919\
        );

    \I__285\ : InMux
    port map (
            O => \N__1925\,
            I => \N__1916\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1922\,
            I => \iterate_regZ0Z_3\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__1919\,
            I => \iterate_regZ0Z_3\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__1916\,
            I => \iterate_regZ0Z_3\
        );

    \I__281\ : IoInMux
    port map (
            O => \N__1909\,
            I => \N__1906\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__1906\,
            I => \N__1903\
        );

    \I__279\ : IoSpan4Mux
    port map (
            O => \N__1903\,
            I => \N__1900\
        );

    \I__278\ : Span4Mux_s0_h
    port map (
            O => \N__1900\,
            I => \N__1897\
        );

    \I__277\ : Span4Mux_h
    port map (
            O => \N__1897\,
            I => \N__1894\
        );

    \I__276\ : Odrv4
    port map (
            O => \N__1894\,
            I => res_out_c_4
        );

    \I__275\ : IoInMux
    port map (
            O => \N__1891\,
            I => \N__1888\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__1888\,
            I => \N__1885\
        );

    \I__273\ : Span4Mux_s2_h
    port map (
            O => \N__1885\,
            I => \N__1882\
        );

    \I__272\ : Span4Mux_v
    port map (
            O => \N__1882\,
            I => \N__1879\
        );

    \I__271\ : Span4Mux_v
    port map (
            O => \N__1879\,
            I => \N__1876\
        );

    \I__270\ : Odrv4
    port map (
            O => \N__1876\,
            I => res_out_c_2
        );

    \I__269\ : IoInMux
    port map (
            O => \N__1873\,
            I => \N__1870\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__1870\,
            I => \N__1867\
        );

    \I__267\ : Span12Mux_s4_h
    port map (
            O => \N__1867\,
            I => \N__1864\
        );

    \I__266\ : Odrv12
    port map (
            O => \N__1864\,
            I => res_out_c_5
        );

    \I__265\ : IoInMux
    port map (
            O => \N__1861\,
            I => \N__1858\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1858\,
            I => \N__1855\
        );

    \I__263\ : Span4Mux_s1_h
    port map (
            O => \N__1855\,
            I => \N__1852\
        );

    \I__262\ : Sp12to4
    port map (
            O => \N__1852\,
            I => \N__1849\
        );

    \I__261\ : Span12Mux_v
    port map (
            O => \N__1849\,
            I => \N__1846\
        );

    \I__260\ : Odrv12
    port map (
            O => \N__1846\,
            I => res_out_c_1
        );

    \I__259\ : CascadeMux
    port map (
            O => \N__1843\,
            I => \N__1840\
        );

    \I__258\ : InMux
    port map (
            O => \N__1840\,
            I => \N__1837\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1837\,
            I => den_reg_i_0
        );

    \I__256\ : InMux
    port map (
            O => \N__1834\,
            I => \N__1831\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1831\,
            I => load_and_iterate_iterate_reg_1_1
        );

    \I__254\ : InMux
    port map (
            O => \N__1828\,
            I => load_and_iterate_iterate_reg_1_cry_0
        );

    \I__253\ : InMux
    port map (
            O => \N__1825\,
            I => \N__1822\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__1822\,
            I => load_and_iterate_iterate_reg_1_2
        );

    \I__251\ : InMux
    port map (
            O => \N__1819\,
            I => load_and_iterate_iterate_reg_1_cry_1
        );

    \I__250\ : IoInMux
    port map (
            O => \N__1816\,
            I => \N__1813\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1813\,
            I => \N__1810\
        );

    \I__248\ : IoSpan4Mux
    port map (
            O => \N__1810\,
            I => \N__1807\
        );

    \I__247\ : Span4Mux_s3_h
    port map (
            O => \N__1807\,
            I => \N__1804\
        );

    \I__246\ : Odrv4
    port map (
            O => \N__1804\,
            I => rmn_out_c_5
        );

    \I__245\ : IoInMux
    port map (
            O => \N__1801\,
            I => \N__1798\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1798\,
            I => \N__1795\
        );

    \I__243\ : IoSpan4Mux
    port map (
            O => \N__1795\,
            I => \N__1792\
        );

    \I__242\ : Span4Mux_s2_h
    port map (
            O => \N__1792\,
            I => \N__1789\
        );

    \I__241\ : Odrv4
    port map (
            O => \N__1789\,
            I => rmn_out_c_6
        );

    \I__240\ : IoInMux
    port map (
            O => \N__1786\,
            I => \N__1783\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__1783\,
            I => \N__1780\
        );

    \I__238\ : IoSpan4Mux
    port map (
            O => \N__1780\,
            I => \N__1777\
        );

    \I__237\ : Span4Mux_s1_h
    port map (
            O => \N__1777\,
            I => \N__1774\
        );

    \I__236\ : Odrv4
    port map (
            O => \N__1774\,
            I => rmn_out_c_0
        );

    \I__235\ : IoInMux
    port map (
            O => \N__1771\,
            I => \N__1768\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__1768\,
            I => \N__1765\
        );

    \I__233\ : Odrv12
    port map (
            O => \N__1765\,
            I => rmn_out_c_2
        );

    \I__232\ : IoInMux
    port map (
            O => \N__1762\,
            I => \N__1759\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__1759\,
            I => \N__1756\
        );

    \I__230\ : IoSpan4Mux
    port map (
            O => \N__1756\,
            I => \N__1753\
        );

    \I__229\ : Span4Mux_s2_h
    port map (
            O => \N__1753\,
            I => \N__1750\
        );

    \I__228\ : Odrv4
    port map (
            O => \N__1750\,
            I => rmn_out_c_1
        );

    \I__227\ : IoInMux
    port map (
            O => \N__1747\,
            I => \N__1744\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1744\,
            I => \N__1741\
        );

    \I__225\ : IoSpan4Mux
    port map (
            O => \N__1741\,
            I => \N__1738\
        );

    \I__224\ : Span4Mux_s3_h
    port map (
            O => \N__1738\,
            I => \N__1735\
        );

    \I__223\ : Span4Mux_v
    port map (
            O => \N__1735\,
            I => \N__1732\
        );

    \I__222\ : Span4Mux_v
    port map (
            O => \N__1732\,
            I => \N__1729\
        );

    \I__221\ : Odrv4
    port map (
            O => \N__1729\,
            I => res_out_c_0
        );

    \I__220\ : IoInMux
    port map (
            O => \N__1726\,
            I => \N__1723\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__1723\,
            I => \N__1720\
        );

    \I__218\ : Span4Mux_s3_h
    port map (
            O => \N__1720\,
            I => \N__1717\
        );

    \I__217\ : Span4Mux_v
    port map (
            O => \N__1717\,
            I => \N__1714\
        );

    \I__216\ : Span4Mux_v
    port map (
            O => \N__1714\,
            I => \N__1711\
        );

    \I__215\ : Odrv4
    port map (
            O => \N__1711\,
            I => res_out_c_3
        );

    \I__214\ : IoInMux
    port map (
            O => \N__1708\,
            I => \N__1705\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__1705\,
            I => \N__1702\
        );

    \I__212\ : Span4Mux_s0_h
    port map (
            O => \N__1702\,
            I => \N__1699\
        );

    \I__211\ : Span4Mux_h
    port map (
            O => \N__1699\,
            I => \N__1696\
        );

    \I__210\ : Odrv4
    port map (
            O => \N__1696\,
            I => res_out_c_7
        );

    \I__209\ : IoInMux
    port map (
            O => \N__1693\,
            I => \N__1690\
        );

    \I__208\ : LocalMux
    port map (
            O => \N__1690\,
            I => \N__1687\
        );

    \I__207\ : Span12Mux_s4_h
    port map (
            O => \N__1687\,
            I => \N__1684\
        );

    \I__206\ : Odrv12
    port map (
            O => \N__1684\,
            I => res_out_c_6
        );

    \I__205\ : InMux
    port map (
            O => \N__1681\,
            I => \N__1678\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__1678\,
            I => \N__1675\
        );

    \I__203\ : Span4Mux_h
    port map (
            O => \N__1675\,
            I => \N__1672\
        );

    \I__202\ : Sp12to4
    port map (
            O => \N__1672\,
            I => \N__1669\
        );

    \I__201\ : Span12Mux_v
    port map (
            O => \N__1669\,
            I => \N__1666\
        );

    \I__200\ : Odrv12
    port map (
            O => \N__1666\,
            I => num_in_c_1
        );

    \I__199\ : InMux
    port map (
            O => \N__1663\,
            I => \N__1660\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1660\,
            I => \N__1657\
        );

    \I__197\ : Span12Mux_v
    port map (
            O => \N__1657\,
            I => \N__1654\
        );

    \I__196\ : Odrv12
    port map (
            O => \N__1654\,
            I => num_in_c_2
        );

    \I__195\ : InMux
    port map (
            O => \N__1651\,
            I => \N__1648\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__1648\,
            I => \N__1645\
        );

    \I__193\ : Span12Mux_s5_h
    port map (
            O => \N__1645\,
            I => \N__1642\
        );

    \I__192\ : Span12Mux_v
    port map (
            O => \N__1642\,
            I => \N__1639\
        );

    \I__191\ : Odrv12
    port map (
            O => \N__1639\,
            I => num_in_c_3
        );

    \I__190\ : InMux
    port map (
            O => \N__1636\,
            I => \N__1633\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__1633\,
            I => \N__1630\
        );

    \I__188\ : Sp12to4
    port map (
            O => \N__1630\,
            I => \N__1627\
        );

    \I__187\ : Span12Mux_v
    port map (
            O => \N__1627\,
            I => \N__1624\
        );

    \I__186\ : Odrv12
    port map (
            O => \N__1624\,
            I => num_in_c_4
        );

    \I__185\ : InMux
    port map (
            O => \N__1621\,
            I => \N__1618\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__1618\,
            I => \N__1615\
        );

    \I__183\ : Span4Mux_h
    port map (
            O => \N__1615\,
            I => \N__1612\
        );

    \I__182\ : Sp12to4
    port map (
            O => \N__1612\,
            I => \N__1609\
        );

    \I__181\ : Span12Mux_v
    port map (
            O => \N__1609\,
            I => \N__1606\
        );

    \I__180\ : Odrv12
    port map (
            O => \N__1606\,
            I => num_in_c_5
        );

    \I__179\ : InMux
    port map (
            O => \N__1603\,
            I => \N__1600\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1600\,
            I => \N__1597\
        );

    \I__177\ : Span4Mux_h
    port map (
            O => \N__1597\,
            I => \N__1594\
        );

    \I__176\ : Sp12to4
    port map (
            O => \N__1594\,
            I => \N__1591\
        );

    \I__175\ : Span12Mux_v
    port map (
            O => \N__1591\,
            I => \N__1588\
        );

    \I__174\ : Odrv12
    port map (
            O => \N__1588\,
            I => num_in_c_6
        );

    \I__173\ : IoInMux
    port map (
            O => \N__1585\,
            I => \N__1582\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1582\,
            I => \N__1579\
        );

    \I__171\ : Span4Mux_s0_h
    port map (
            O => \N__1579\,
            I => \N__1576\
        );

    \I__170\ : Span4Mux_v
    port map (
            O => \N__1576\,
            I => \N__1573\
        );

    \I__169\ : Span4Mux_h
    port map (
            O => \N__1573\,
            I => \N__1570\
        );

    \I__168\ : Odrv4
    port map (
            O => \N__1570\,
            I => rmn_out_c_7
        );

    \I__167\ : IoInMux
    port map (
            O => \N__1567\,
            I => \N__1564\
        );

    \I__166\ : LocalMux
    port map (
            O => \N__1564\,
            I => \N__1561\
        );

    \I__165\ : Odrv12
    port map (
            O => \N__1561\,
            I => rmn_out_c_3
        );

    \I__164\ : IoInMux
    port map (
            O => \N__1558\,
            I => \N__1555\
        );

    \I__163\ : LocalMux
    port map (
            O => \N__1555\,
            I => \N__1552\
        );

    \I__162\ : Span4Mux_s0_h
    port map (
            O => \N__1552\,
            I => \N__1549\
        );

    \I__161\ : Span4Mux_h
    port map (
            O => \N__1549\,
            I => \N__1546\
        );

    \I__160\ : Odrv4
    port map (
            O => \N__1546\,
            I => rmn_out_c_4
        );

    \I__159\ : InMux
    port map (
            O => \N__1543\,
            I => \N__1540\
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1540\,
            I => \N__1537\
        );

    \I__157\ : Sp12to4
    port map (
            O => \N__1537\,
            I => \N__1534\
        );

    \I__156\ : Span12Mux_v
    port map (
            O => \N__1534\,
            I => \N__1531\
        );

    \I__155\ : Odrv12
    port map (
            O => \N__1531\,
            I => rst_in_n_c
        );

    \I__154\ : IoInMux
    port map (
            O => \N__1528\,
            I => \N__1525\
        );

    \I__153\ : LocalMux
    port map (
            O => \N__1525\,
            I => \N__1522\
        );

    \I__152\ : Span4Mux_s3_h
    port map (
            O => \N__1522\,
            I => \N__1519\
        );

    \I__151\ : Span4Mux_v
    port map (
            O => \N__1519\,
            I => \N__1516\
        );

    \I__150\ : Odrv4
    port map (
            O => \N__1516\,
            I => rst_in_n_c_i
        );

    \I__149\ : InMux
    port map (
            O => \N__1513\,
            I => \N__1510\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__1510\,
            I => \N__1507\
        );

    \I__147\ : Span12Mux_h
    port map (
            O => \N__1507\,
            I => \N__1504\
        );

    \I__146\ : Span12Mux_v
    port map (
            O => \N__1504\,
            I => \N__1501\
        );

    \I__145\ : Odrv12
    port map (
            O => \N__1501\,
            I => den_in_c_0
        );

    \I__144\ : InMux
    port map (
            O => \N__1498\,
            I => \N__1495\
        );

    \I__143\ : LocalMux
    port map (
            O => \N__1495\,
            I => \N__1492\
        );

    \I__142\ : Sp12to4
    port map (
            O => \N__1492\,
            I => \N__1489\
        );

    \I__141\ : Span12Mux_v
    port map (
            O => \N__1489\,
            I => \N__1486\
        );

    \I__140\ : Odrv12
    port map (
            O => \N__1486\,
            I => den_in_c_5
        );

    \I__139\ : InMux
    port map (
            O => \N__1483\,
            I => \N__1480\
        );

    \I__138\ : LocalMux
    port map (
            O => \N__1480\,
            I => \N__1477\
        );

    \I__137\ : Span4Mux_v
    port map (
            O => \N__1477\,
            I => \N__1474\
        );

    \I__136\ : Span4Mux_h
    port map (
            O => \N__1474\,
            I => \N__1471\
        );

    \I__135\ : Span4Mux_v
    port map (
            O => \N__1471\,
            I => \N__1468\
        );

    \I__134\ : Span4Mux_v
    port map (
            O => \N__1468\,
            I => \N__1465\
        );

    \I__133\ : Odrv4
    port map (
            O => \N__1465\,
            I => den_in_c_6
        );

    \I__132\ : CascadeMux
    port map (
            O => \N__1462\,
            I => \N__1459\
        );

    \I__131\ : InMux
    port map (
            O => \N__1459\,
            I => \N__1456\
        );

    \I__130\ : LocalMux
    port map (
            O => \N__1456\,
            I => \N__1453\
        );

    \I__129\ : Span4Mux_h
    port map (
            O => \N__1453\,
            I => \N__1450\
        );

    \I__128\ : Sp12to4
    port map (
            O => \N__1450\,
            I => \N__1447\
        );

    \I__127\ : Span12Mux_v
    port map (
            O => \N__1447\,
            I => \N__1444\
        );

    \I__126\ : Odrv12
    port map (
            O => \N__1444\,
            I => num_in_c_0
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => iterate_ena_li,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_13_0_\
        );

    \rst_in_n_ibuf_RNI1DMA_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__1528\,
            GLOBALBUFFEROUTPUT => rst_in_n_c_i_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \rst_in_n_ibuf_RNI1DMA_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__1543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rst_in_n_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \den_reg_0_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1513\,
            lcout => \den_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2790\,
            ce => \N__2891\,
            sr => \N__2756\
        );

    \den_reg_5_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1498\,
            lcout => \den_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2790\,
            ce => \N__2891\,
            sr => \N__2756\
        );

    \den_reg_6_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1483\,
            lcout => \den_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2790\,
            ce => \N__2891\,
            sr => \N__2756\
        );

    \iterate_reg_0_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__2895\,
            in1 => \N__2576\,
            in2 => \N__1462\,
            in3 => \N__2013\,
            lcout => \iterate_regZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2789\,
            ce => \N__2472\,
            sr => \N__2758\
        );

    \iterate_reg_1_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__1681\,
            in1 => \N__2896\,
            in2 => \_gnd_net_\,
            in3 => \N__1834\,
            lcout => \iterate_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2789\,
            ce => \N__2472\,
            sr => \N__2758\
        );

    \iterate_reg_2_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__2892\,
            in1 => \N__1663\,
            in2 => \_gnd_net_\,
            in3 => \N__1825\,
            lcout => \iterate_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2789\,
            ce => \N__2472\,
            sr => \N__2758\
        );

    \iterate_reg_3_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__1651\,
            in1 => \N__2897\,
            in2 => \_gnd_net_\,
            in3 => \N__2098\,
            lcout => \iterate_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2789\,
            ce => \N__2472\,
            sr => \N__2758\
        );

    \iterate_reg_4_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__2893\,
            in1 => \N__1636\,
            in2 => \_gnd_net_\,
            in3 => \N__2089\,
            lcout => \iterate_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2789\,
            ce => \N__2472\,
            sr => \N__2758\
        );

    \iterate_reg_5_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__1621\,
            in1 => \N__2898\,
            in2 => \_gnd_net_\,
            in3 => \N__2071\,
            lcout => \iterate_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2789\,
            ce => \N__2472\,
            sr => \N__2758\
        );

    \iterate_reg_6_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__2894\,
            in1 => \N__1603\,
            in2 => \_gnd_net_\,
            in3 => \N__2053\,
            lcout => \iterate_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2789\,
            ce => \N__2472\,
            sr => \N__2758\
        );

    \rmn_outZ0Z_7_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2446\,
            lcout => rmn_out_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => \N__2631\,
            sr => \N__2759\
        );

    \rmn_outZ0Z_3_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1927\,
            lcout => rmn_out_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => \N__2631\,
            sr => \N__2759\
        );

    \rmn_outZ0Z_4_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2196\,
            lcout => rmn_out_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => \N__2631\,
            sr => \N__2759\
        );

    \rmn_outZ0Z_5_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2167\,
            lcout => rmn_out_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => \N__2631\,
            sr => \N__2759\
        );

    \rmn_outZ0Z_6_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2140\,
            lcout => rmn_out_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => \N__2631\,
            sr => \N__2759\
        );

    \rmn_outZ0Z_0_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2014\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => rmn_out_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => \N__2631\,
            sr => \N__2759\
        );

    \rmn_outZ0Z_2_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1954\,
            lcout => rmn_out_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => \N__2631\,
            sr => \N__2759\
        );

    \rmn_outZ0Z_1_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1981\,
            lcout => rmn_out_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2791\,
            ce => \N__2631\,
            sr => \N__2759\
        );

    \res_outZ0Z_0_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2281\,
            lcout => res_out_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2632\,
            sr => \N__2760\
        );

    \res_outZ0Z_3_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2236\,
            lcout => res_out_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2632\,
            sr => \N__2760\
        );

    \res_outZ0Z_7_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2485\,
            lcout => res_out_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2632\,
            sr => \N__2760\
        );

    \res_outZ0Z_6_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2503\,
            lcout => res_out_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2632\,
            sr => \N__2760\
        );

    \res_outZ0Z_4_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2221\,
            lcout => res_out_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2632\,
            sr => \N__2760\
        );

    \res_outZ0Z_2_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2251\,
            lcout => res_out_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2632\,
            sr => \N__2760\
        );

    \res_outZ0Z_5_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2518\,
            lcout => res_out_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2632\,
            sr => \N__2760\
        );

    \res_outZ0Z_1_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2266\,
            lcout => res_out_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2793\,
            ce => \N__2632\,
            sr => \N__2760\
        );

    \den_reg_sbtinv_5_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2344\,
            lcout => den_reg_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \den_reg_sbtinv_6_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2310\,
            lcout => den_reg_i_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \load_and_iterate_iterate_reg_1_cry_0_c_inv_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2569\,
            in1 => \N__2012\,
            in2 => \N__1843\,
            in3 => \_gnd_net_\,
            lcout => den_reg_i_0,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => load_and_iterate_iterate_reg_1_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \iterate_reg_RNO_0_1_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1980\,
            in2 => \N__2404\,
            in3 => \N__1828\,
            lcout => load_and_iterate_iterate_reg_1_1,
            ltout => OPEN,
            carryin => load_and_iterate_iterate_reg_1_cry_0,
            carryout => load_and_iterate_iterate_reg_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \iterate_reg_RNO_0_2_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1953\,
            in2 => \N__2395\,
            in3 => \N__1819\,
            lcout => load_and_iterate_iterate_reg_1_2,
            ltout => OPEN,
            carryin => load_and_iterate_iterate_reg_1_cry_1,
            carryout => load_and_iterate_iterate_reg_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \iterate_reg_RNO_0_3_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1926\,
            in2 => \N__2419\,
            in3 => \N__2092\,
            lcout => load_and_iterate_iterate_reg_1_3,
            ltout => OPEN,
            carryin => load_and_iterate_iterate_reg_1_cry_2,
            carryout => load_and_iterate_iterate_reg_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \iterate_reg_RNO_0_4_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2410\,
            in2 => \N__2197\,
            in3 => \N__2083\,
            lcout => load_and_iterate_iterate_reg_1_4,
            ltout => OPEN,
            carryin => load_and_iterate_iterate_reg_1_cry_3,
            carryout => load_and_iterate_iterate_reg_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \iterate_reg_RNO_0_5_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2166\,
            in2 => \N__2080\,
            in3 => \N__2065\,
            lcout => load_and_iterate_iterate_reg_1_5,
            ltout => OPEN,
            carryin => load_and_iterate_iterate_reg_1_cry_4,
            carryout => load_and_iterate_iterate_reg_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \iterate_reg_RNO_0_6_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2139\,
            in2 => \N__2062\,
            in3 => \N__2047\,
            lcout => load_and_iterate_iterate_reg_1_6,
            ltout => OPEN,
            carryin => load_and_iterate_iterate_reg_1_cry_5,
            carryout => load_and_iterate_iterate_reg_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \iterate_reg_7_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__2890\,
            in1 => \N__2425\,
            in2 => \N__2044\,
            in3 => \N__2017\,
            lcout => \iterate_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2794\,
            ce => \N__2473\,
            sr => \N__2757\
        );

    \is_higher_than_un1_iterate_reg_cry_0_c_inv_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2568\,
            in2 => \N__1990\,
            in3 => \N__2011\,
            lcout => iterate_reg_i_0,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => is_higher_than_un1_iterate_reg_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \is_higher_than_un1_iterate_reg_cry_1_c_inv_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2611\,
            in2 => \N__1963\,
            in3 => \N__1979\,
            lcout => iterate_reg_i_1,
            ltout => OPEN,
            carryin => is_higher_than_un1_iterate_reg_cry_0,
            carryout => is_higher_than_un1_iterate_reg_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \is_higher_than_un1_iterate_reg_cry_2_c_inv_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3070\,
            in2 => \N__1936\,
            in3 => \N__1952\,
            lcout => iterate_reg_i_2,
            ltout => OPEN,
            carryin => is_higher_than_un1_iterate_reg_cry_1,
            carryout => is_higher_than_un1_iterate_reg_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \is_higher_than_un1_iterate_reg_cry_3_c_inv_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3107\,
            in2 => \N__2206\,
            in3 => \N__1925\,
            lcout => iterate_reg_i_3,
            ltout => OPEN,
            carryin => is_higher_than_un1_iterate_reg_cry_2,
            carryout => is_higher_than_un1_iterate_reg_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \is_higher_than_un1_iterate_reg_cry_4_c_inv_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2650\,
            in2 => \N__2176\,
            in3 => \N__2192\,
            lcout => iterate_reg_i_4,
            ltout => OPEN,
            carryin => is_higher_than_un1_iterate_reg_cry_3,
            carryout => is_higher_than_un1_iterate_reg_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \is_higher_than_un1_iterate_reg_cry_5_c_inv_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2345\,
            in2 => \N__2149\,
            in3 => \N__2165\,
            lcout => iterate_reg_i_5,
            ltout => OPEN,
            carryin => is_higher_than_un1_iterate_reg_cry_4,
            carryout => is_higher_than_un1_iterate_reg_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \is_higher_than_un1_iterate_reg_cry_6_c_inv_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2309\,
            in2 => \N__2122\,
            in3 => \N__2138\,
            lcout => iterate_reg_i_6,
            ltout => OPEN,
            carryin => is_higher_than_un1_iterate_reg_cry_5,
            carryout => is_higher_than_un1_iterate_reg_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \is_higher_than_un1_iterate_reg_cry_7_c_inv_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2368\,
            in2 => \N__2113\,
            in3 => \N__2441\,
            lcout => iterate_reg_i_7,
            ltout => OPEN,
            carryin => is_higher_than_un1_iterate_reg_cry_6,
            carryout => iterate_ena_li,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \iterate_ena_li_THRU_LUT4_0_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2104\,
            lcout => \iterate_ena_li_THRU_CO\,
            ltout => \iterate_ena_li_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_state_RNO_0_3_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2985\,
            in2 => \N__2101\,
            in3 => \N__2922\,
            lcout => current_state_ns_i_rn_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \is_higher_than_un1_iterate_reg_cry_7_c_RNIREHR_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2989\,
            in2 => \_gnd_net_\,
            in3 => \N__2289\,
            lcout => \N_4_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_state_RNO_1_3_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__2923\,
            in1 => \N__2370\,
            in2 => \N__2998\,
            in3 => \N__2322\,
            lcout => current_state_ns_i_sn_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_state_RNO_3_3_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2613\,
            in1 => \N__3075\,
            in2 => \N__3109\,
            in3 => \N__2577\,
            lcout => is_den_zero_un5_den_reg_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_state_RNO_2_3_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__2653\,
            in1 => \N__2346\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => is_den_zero_un5_den_reg_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_state_RNO_1_2_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2371\,
            in1 => \N__2652\,
            in2 => \N__2350\,
            in3 => \N__2323\,
            lcout => o2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \is_higher_than_un1_iterate_reg_cry_7_c_RNI6DU81_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2864\,
            in2 => \N__2293\,
            in3 => \N__2984\,
            lcout => counter_cnte_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_cnt_0_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2863\,
            in1 => \N__2280\,
            in2 => \_gnd_net_\,
            in3 => \N__2269\,
            lcout => \counter_cntZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => counter_cnt_cry_0,
            clk => \N__2795\,
            ce => \N__2468\,
            sr => \N__2762\
        );

    \counter_cnt_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2856\,
            in1 => \N__2265\,
            in2 => \_gnd_net_\,
            in3 => \N__2254\,
            lcout => \counter_cntZ0Z_1\,
            ltout => OPEN,
            carryin => counter_cnt_cry_0,
            carryout => counter_cnt_cry_1,
            clk => \N__2795\,
            ce => \N__2468\,
            sr => \N__2762\
        );

    \counter_cnt_2_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2859\,
            in1 => \N__2250\,
            in2 => \_gnd_net_\,
            in3 => \N__2239\,
            lcout => \counter_cntZ0Z_2\,
            ltout => OPEN,
            carryin => counter_cnt_cry_1,
            carryout => counter_cnt_cry_2,
            clk => \N__2795\,
            ce => \N__2468\,
            sr => \N__2762\
        );

    \counter_cnt_3_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2857\,
            in1 => \N__2235\,
            in2 => \_gnd_net_\,
            in3 => \N__2224\,
            lcout => \counter_cntZ0Z_3\,
            ltout => OPEN,
            carryin => counter_cnt_cry_2,
            carryout => counter_cnt_cry_3,
            clk => \N__2795\,
            ce => \N__2468\,
            sr => \N__2762\
        );

    \counter_cnt_4_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2860\,
            in1 => \N__2220\,
            in2 => \_gnd_net_\,
            in3 => \N__2209\,
            lcout => \counter_cntZ0Z_4\,
            ltout => OPEN,
            carryin => counter_cnt_cry_3,
            carryout => counter_cnt_cry_4,
            clk => \N__2795\,
            ce => \N__2468\,
            sr => \N__2762\
        );

    \counter_cnt_5_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2858\,
            in1 => \N__2517\,
            in2 => \_gnd_net_\,
            in3 => \N__2506\,
            lcout => \counter_cntZ0Z_5\,
            ltout => OPEN,
            carryin => counter_cnt_cry_4,
            carryout => counter_cnt_cry_5,
            clk => \N__2795\,
            ce => \N__2468\,
            sr => \N__2762\
        );

    \counter_cnt_6_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2861\,
            in1 => \N__2502\,
            in2 => \_gnd_net_\,
            in3 => \N__2491\,
            lcout => \counter_cntZ0Z_6\,
            ltout => OPEN,
            carryin => counter_cnt_cry_5,
            carryout => counter_cnt_cry_6,
            clk => \N__2795\,
            ce => \N__2468\,
            sr => \N__2762\
        );

    \counter_cnt_7_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__2484\,
            in1 => \N__2862\,
            in2 => \_gnd_net_\,
            in3 => \N__2488\,
            lcout => \counter_cntZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2795\,
            ce => \N__2468\,
            sr => \N__2762\
        );

    \iterate_reg_RNO_0_7_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2369\,
            in2 => \_gnd_net_\,
            in3 => \N__2442\,
            lcout => load_and_iterate_iterate_reg_1_axb_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \den_reg_sbtinv_3_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3100\,
            lcout => den_reg_i_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \den_reg_sbtinv_4_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2651\,
            lcout => den_reg_i_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \den_reg_sbtinv_1_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2612\,
            lcout => den_reg_i_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \den_reg_sbtinv_2_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3071\,
            lcout => den_reg_i_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \den_reg_7_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2386\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \den_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2792\,
            ce => \N__2899\,
            sr => \N__2761\
        );

    \den_reg_2_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \den_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2792\,
            ce => \N__2899\,
            sr => \N__2761\
        );

    \den_reg_1_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2710\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \den_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2792\,
            ce => \N__2899\,
            sr => \N__2761\
        );

    \den_reg_3_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2689\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \den_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2792\,
            ce => \N__2899\,
            sr => \N__2761\
        );

    \den_reg_4_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2668\,
            lcout => \den_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2792\,
            ce => \N__2899\,
            sr => \N__2761\
        );

    \current_state_4_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2630\,
            lcout => \resultOk_out_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2796\,
            ce => 'H',
            sr => \N__2763\
        );

    \current_state_2_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3049\,
            in1 => \N__2614\,
            in2 => \N__2590\,
            in3 => \N__2581\,
            lcout => \divZero_out_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2796\,
            ce => 'H',
            sr => \N__2763\
        );

    \current_state_3_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111001011111010"
        )
    port map (
            in0 => \N__2545\,
            in1 => \N__2539\,
            in2 => \N__2533\,
            in3 => \N__2524\,
            lcout => \current_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2796\,
            ce => 'H',
            sr => \N__2763\
        );

    \current_state_1_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2871\,
            lcout => \current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2796\,
            ce => 'H',
            sr => \N__2763\
        );

    \current_state_RNO_0_5_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__3015\,
            in1 => \N__2962\,
            in2 => \N__3150\,
            in3 => \N__3120\,
            lcout => current_state_ns_i_0_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_state_RNO_0_2_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__2924\,
            in1 => \N__3108\,
            in2 => \_gnd_net_\,
            in3 => \N__3076\,
            lcout => m4_e_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \running_out_obuf_RNO_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__2925\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3003\,
            lcout => \N_58_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_state_5_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__2932\,
            in1 => \N__3025\,
            in2 => \N__3004\,
            in3 => \N__2957\,
            lcout => \current_stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2797\,
            ce => 'H',
            sr => \N__2764\
        );

    \current_state_0_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__3016\,
            in1 => \N__2999\,
            in2 => \N__2961\,
            in3 => \N__2931\,
            lcout => \current_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2797\,
            ce => 'H',
            sr => \N__2764\
        );
end \INTERFACE\;
