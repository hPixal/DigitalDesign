library ieee;
use ieee.std_logic_1164.all; 

entity Valvula is
    port(
        act_valvula : in std_logic
        );
end entity;
