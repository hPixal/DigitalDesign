library ieee;
use ieee.std_logic_1164.all;

entity Bomba is
port(
    act_bomba : in std_logic
);
end entity;