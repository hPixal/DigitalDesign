package parametersPackage is
    constant NCOBITS : integer :=  4;
    constant FREQCONTROLBITS : integer := 3;
end parametersPackage;
