library ieee;
use ieee.std_logic_1164.all;
---use ieee.std_logic_arth.all;
---use ieee.std_logic_unsigned.all;

entity tipoJK_tb is
end entity;

architecture tipoJK_tb of tipoJK_tb is
    component tipoJK